library IEEE;
USE ieee.std_logic_1164.all;

ENTITY StateMachine is
PORT (
      clock : 	IN STD_LOGIC;
      reset : 	IN STD_LOGIC;
      inbus :	IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      outbus :	OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ENTITY;

-- Architecture definition for the SimpleFSM entity
Architecture behave of StateMachine is
TYPE State_type IS (INIT, TEST1, ADD, SUB, Q0, TEST_COUNT7, SHIFT, TEST2, OUTPUT, STOP);  -- Define the states
	SIGNAL State : State_Type;    -- Create a signal that uses the different states
	SIGNAL A,Q,M: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL count7: STD_LOGIC;
	
-- Component declarations region				    
COMPONENT adder IS
	PORT(clock, c_in: IN STD_LOGIC;
		x,y: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		z: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		c_out: OUT STD_LOGIC);
END COMPONENT;

COMPONENT shiftRegister IS
	GENERIC( n: INTEGER);
	PORT(clock: IN STD_LOGIC;
		intrare: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		iesire: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0));
END COMPONENT;

COMPONENT controlUnit IS
	PORT(clock, begin_sgn, q0, count7: IN BIT;
		end_sgn,c0,c1,c2,c3,c4,c5,c6,c7,c8: OUT BIT);
END COMPONENT;

COMPONENT counter IS
	PORT(clock: IN STD_LOGIC;
		in_val: IN INTEGER;
		out_val: OUT INTEGER;
		count7: OUT STD_LOGIC);
END COMPONENT;

	SIGNAL s: STD_LOGIC;
	SIGNAL sum_out, compl2 : std_logic_vector(7 downto 0);
	SIGNAL shift_in, shift_out : std_logic_vector(15 downto 0);
-- end region

BEGIN 
-- Component instantiation
shiftReg: shiftRegister 
	generic map ( n => 16 )
	port map (clock => clock,
		intrare => shift_in,
		iesire => shift_out);

adder_entity: adder 
	port map(clock => clock, 
		c_in => '0',
		x => a,
		y => m,
		z => a,
		c_out => s);

subtractor_entity: adder 
	port map(clock => clock, 
		c_in => '0',
		x => a,
		y => compl2,
		z => a,
		c_out => s);
--end region


  PROCESS (clock, reset) 
	VARIABLE c0,c1,c2,c3,c4,c5,c6,c7,c8,at_end: STD_LOGIC := '0';
	VARIABLE count: INTEGER;

  BEGIN 
    IF (reset = '1') THEN            -- upon reset, set the state to INIT
    	State <= INIT;
 
    ELSIF rising_edge(clock) THEN   

		CASE State IS

			WHEN INIT => 
				at_end:='0';
				s<='0';
				count:=0;

				A<=inbus(15 downto 8);
				Q(7 downto 1)<=inbus(7 downto 1);
				Q(0)<='0';
				M<=inbus(7 downto 0);
				State<=TEST1;

			WHEN TEST1 => 
				IF s='1' THEN 
					State <= ADD; 
				ELSE
					State <= SUB;
				END IF; 

			WHEN ADD => 
				--add				
				
				IF (at_end = '1') THEN
					State <= OUTPUT;
				ELSE
					State <=Q0;
				END IF; 

			WHEN SUB => 
				compl2 <= m;
				-- sub
				State <= Q0; 

			WHEN Q0 => 
				Q(0) <= NOT(s); 

			WHEN TEST_COUNT7 => 
				IF count7='1' THEN 
					State <= SHIFT; 
				ELSE 
					State <= TEST2; 
				END IF; 

			WHEN SHIFT => 
				shift_in(15 downto 8)<=a;
				shift_in(7 downto 0)<=q;

				--shifting
				
				s<=shift_out(15);
				a<=shift_out(14 downto 7);
				q(7 downto 1)<=shift_out(6 downto 0);
				q(0) <= '0';
				count:=count+1;
				if(count = 7) then count7<='1'; end if;

			WHEN TEST2 => 
				IF s='1' THEN 
					at_end:='1';
					State <= ADD; 
				ELSE 
					State <= OUTPUT; 
				END IF; 
			
			WHEN OUTPUT => 
				Outbus(15 downto 8) <= Q;
				Outbus(7 downto 0) <= A;
				State <= STOP; 
				
			WHEN STOP =>

			WHEN others =>
				State <= INIT;
		END CASE; 
    END IF; 
  END PROCESS;
  
END behave;
